//////////////
//conf_1
assign I_configs[0][1] = I_in_temp[0];
assign I_configs[1][1] = I_in_temp[1];
assign I_configs[2][1] = I_in_temp[2];
assign I_configs[3][1] = I_in_temp[3];
assign I_configs[4][1] = I_in_temp[4];
assign I_configs[5][1] = I_in_temp[5];
assign I_configs[6][1] = I_in_temp[6];
assign I_configs[7][1] = I_in_temp[7];
assign I_configs[8][1] = I_in_temp[0];
assign I_configs[9][1] = I_in_temp[1];
assign I_configs[10][1] = I_in_temp[2];
assign I_configs[11][1] = I_in_temp[3];
assign I_configs[12][1] = I_in_temp[4];
assign I_configs[13][1] = I_in_temp[5];
assign I_configs[14][1] = I_in_temp[6];
assign I_configs[15][1] = I_in_temp[7];
assign I_configs[16][1] = I_in_temp[0];
assign I_configs[17][1] = I_in_temp[1];
assign I_configs[18][1] = I_in_temp[2];
assign I_configs[19][1] = I_in_temp[3];
assign I_configs[20][1] = I_in_temp[4];
assign I_configs[21][1] = I_in_temp[5];
assign I_configs[22][1] = I_in_temp[6];
assign I_configs[23][1] = I_in_temp[7];
assign I_configs[24][1] = I_in_temp[0];
assign I_configs[25][1] = I_in_temp[1];
assign I_configs[26][1] = I_in_temp[2];
assign I_configs[27][1] = I_in_temp[3];
assign I_configs[28][1] = I_in_temp[4];
assign I_configs[29][1] = I_in_temp[5];
assign I_configs[30][1] = I_in_temp[6];
assign I_configs[31][1] = I_in_temp[7];
assign Res_configs[0][1] = Res_cas_in_temp[0];
assign Res_configs[1][1] = Res_cascade[0];
assign Res_configs[2][1] = Res_cascade[1];
assign Res_configs[3][1] = Res_cascade[2];
assign Res_configs[4][1] = Res_cas_in_temp[1];
assign Res_configs[5][1] = Res_cascade[4];
assign Res_configs[6][1] = Res_cascade[5];
assign Res_configs[7][1] = Res_cascade[6];
assign Res_configs[8][1] = Res_cas_in_temp[2];
assign Res_configs[9][1] = Res_cascade[8];
assign Res_configs[10][1] = Res_cascade[9];
assign Res_configs[11][1] = Res_cascade[10];
assign Res_configs[12][1] = Res_cas_in_temp[3];
assign Res_configs[13][1] = Res_cascade[12];
assign Res_configs[14][1] = Res_cascade[13];
assign Res_configs[15][1] = Res_cascade[14];
assign Res_configs[16][1] = Res_cas_in_temp[4];
assign Res_configs[17][1] = Res_cascade[16];
assign Res_configs[18][1] = Res_cascade[17];
assign Res_configs[19][1] = Res_cascade[18];
assign Res_configs[20][1] = Res_cas_in_temp[5];
assign Res_configs[21][1] = Res_cascade[20];
assign Res_configs[22][1] = Res_cascade[21];
assign Res_configs[23][1] = Res_cascade[22];
assign Res_configs[24][1] = Res_cas_in_temp[6];
assign Res_configs[25][1] = Res_cascade[24];
assign Res_configs[26][1] = Res_cascade[25];
assign Res_configs[27][1] = Res_cascade[26];
assign Res_configs[28][1] = Res_cas_in_temp[7];
assign Res_configs[29][1] = Res_cascade[28];
assign Res_configs[30][1] = Res_cascade[29];
assign Res_configs[31][1] = Res_cascade[30];
assign Res_out_temp[0][1] = {RES_W{1'bx}};
assign Res_out_temp[1][1] = Res_cascade[4];
assign Res_out_temp[2][1] = {RES_W{1'bx}};
assign Res_out_temp[3][1] = Res_cascade[8];
assign Res_out_temp[4][1] = {RES_W{1'bx}};
assign Res_out_temp[5][1] = Res_cascade[12];
assign Res_out_temp[6][1] = {RES_W{1'bx}};
assign Res_out_temp[7][1] = Res_cascade[16];
assign Res_out_temp[8][1] = {RES_W{1'bx}};
assign Res_out_temp[9][1] = Res_cascade[20];
assign Res_out_temp[10][1] = {RES_W{1'bx}};
assign Res_out_temp[11][1] = Res_cascade[24];
assign Res_out_temp[12][1] = {RES_W{1'bx}};
assign Res_out_temp[13][1] = Res_cascade[28];
assign Res_out_temp[14][1] = {RES_W{1'bx}};
assign Res_out_temp[15][1] = Res_cascade[32];
//////////////
//conf_0
assign I_configs[0][0] = I_in_temp[0];
assign I_configs[1][0] = I_cascade[0];
assign I_configs[2][0] = I_in_temp[1];
assign I_configs[3][0] = I_cascade[2];
assign I_configs[4][0] = I_in_temp[2];
assign I_configs[5][0] = I_cascade[4];
assign I_configs[6][0] = I_in_temp[3];
assign I_configs[7][0] = I_cascade[6];
assign I_configs[8][0] = I_in_temp[0];
assign I_configs[9][0] = I_cascade[8];
assign I_configs[10][0] = I_in_temp[1];
assign I_configs[11][0] = I_cascade[10];
assign I_configs[12][0] = I_in_temp[2];
assign I_configs[13][0] = I_cascade[12];
assign I_configs[14][0] = I_in_temp[3];
assign I_configs[15][0] = I_cascade[14];
assign I_configs[16][0] = I_in_temp[0];
assign I_configs[17][0] = I_cascade[16];
assign I_configs[18][0] = I_in_temp[1];
assign I_configs[19][0] = I_cascade[18];
assign I_configs[20][0] = I_in_temp[2];
assign I_configs[21][0] = I_cascade[20];
assign I_configs[22][0] = I_in_temp[3];
assign I_configs[23][0] = I_cascade[22];
assign I_configs[24][0] = I_in_temp[0];
assign I_configs[25][0] = I_cascade[24];
assign I_configs[26][0] = I_in_temp[1];
assign I_configs[27][0] = I_cascade[26];
assign I_configs[28][0] = I_in_temp[2];
assign I_configs[29][0] = I_cascade[28];
assign I_configs[30][0] = I_in_temp[3];
assign I_configs[31][0] = I_cascade[30];
assign Res_configs[0][0] = Res_cas_in_temp[0];
assign Res_configs[1][0] = Res_cascade[0];
assign Res_configs[2][0] = Res_cascade[1];
assign Res_configs[3][0] = Res_cascade[2];
assign Res_configs[4][0] = Res_cas_in_temp[1];
assign Res_configs[5][0] = Res_cascade[4];
assign Res_configs[6][0] = Res_cascade[5];
assign Res_configs[7][0] = Res_cascade[6];
assign Res_configs[8][0] = Res_cas_in_temp[2];
assign Res_configs[9][0] = Res_cascade[8];
assign Res_configs[10][0] = Res_cascade[9];
assign Res_configs[11][0] = Res_cascade[10];
assign Res_configs[12][0] = Res_cas_in_temp[3];
assign Res_configs[13][0] = Res_cascade[12];
assign Res_configs[14][0] = Res_cascade[13];
assign Res_configs[15][0] = Res_cascade[14];
assign Res_configs[16][0] = Res_cas_in_temp[4];
assign Res_configs[17][0] = Res_cascade[16];
assign Res_configs[18][0] = Res_cascade[17];
assign Res_configs[19][0] = Res_cascade[18];
assign Res_configs[20][0] = Res_cas_in_temp[5];
assign Res_configs[21][0] = Res_cascade[20];
assign Res_configs[22][0] = Res_cascade[21];
assign Res_configs[23][0] = Res_cascade[22];
assign Res_configs[24][0] = Res_cas_in_temp[6];
assign Res_configs[25][0] = Res_cascade[24];
assign Res_configs[26][0] = Res_cascade[25];
assign Res_configs[27][0] = Res_cascade[26];
assign Res_configs[28][0] = Res_cas_in_temp[7];
assign Res_configs[29][0] = Res_cascade[28];
assign Res_configs[30][0] = Res_cascade[29];
assign Res_configs[31][0] = Res_cascade[30];
assign Res_out_temp[0][0] = {RES_W{1'bx}};
assign Res_out_temp[1][0] = Res_cascade[4];
assign Res_out_temp[2][0] = {RES_W{1'bx}};
assign Res_out_temp[3][0] = Res_cascade[8];
assign Res_out_temp[4][0] = {RES_W{1'bx}};
assign Res_out_temp[5][0] = Res_cascade[12];
assign Res_out_temp[6][0] = {RES_W{1'bx}};
assign Res_out_temp[7][0] = Res_cascade[16];
assign Res_out_temp[8][0] = {RES_W{1'bx}};
assign Res_out_temp[9][0] = Res_cascade[20];
assign Res_out_temp[10][0] = {RES_W{1'bx}};
assign Res_out_temp[11][0] = Res_cascade[24];
assign Res_out_temp[12][0] = {RES_W{1'bx}};
assign Res_out_temp[13][0] = Res_cascade[28];
assign Res_out_temp[14][0] = {RES_W{1'bx}};
assign Res_out_temp[15][0] = Res_cascade[32];
//////////////
//conf_3
assign I_configs[0][3] = I_in_temp[0];
assign I_configs[1][3] = I_in_temp[1];
assign I_configs[2][3] = I_in_temp[2];
assign I_configs[3][3] = I_in_temp[3];
assign I_configs[4][3] = I_in_temp[4];
assign I_configs[5][3] = I_in_temp[5];
assign I_configs[6][3] = I_in_temp[6];
assign I_configs[7][3] = I_in_temp[7];
assign I_configs[8][3] = I_in_temp[0];
assign I_configs[9][3] = I_in_temp[1];
assign I_configs[10][3] = I_in_temp[2];
assign I_configs[11][3] = I_in_temp[3];
assign I_configs[12][3] = I_in_temp[4];
assign I_configs[13][3] = I_in_temp[5];
assign I_configs[14][3] = I_in_temp[6];
assign I_configs[15][3] = I_in_temp[7];
assign I_configs[16][3] = I_in_temp[0];
assign I_configs[17][3] = I_in_temp[1];
assign I_configs[18][3] = I_in_temp[2];
assign I_configs[19][3] = I_in_temp[3];
assign I_configs[20][3] = I_in_temp[4];
assign I_configs[21][3] = I_in_temp[5];
assign I_configs[22][3] = I_in_temp[6];
assign I_configs[23][3] = I_in_temp[7];
assign I_configs[24][3] = I_in_temp[0];
assign I_configs[25][3] = I_in_temp[1];
assign I_configs[26][3] = I_in_temp[2];
assign I_configs[27][3] = I_in_temp[3];
assign I_configs[28][3] = I_in_temp[4];
assign I_configs[29][3] = I_in_temp[5];
assign I_configs[30][3] = I_in_temp[6];
assign I_configs[31][3] = I_in_temp[7];
assign Res_configs[0][3] = Res_cas_in_temp[0];
assign Res_configs[1][3] = Res_cascade[0];
assign Res_configs[2][3] = Res_cas_in_temp[1];
assign Res_configs[3][3] = Res_cascade[2];
assign Res_configs[4][3] = Res_cas_in_temp[2];
assign Res_configs[5][3] = Res_cascade[4];
assign Res_configs[6][3] = Res_cas_in_temp[3];
assign Res_configs[7][3] = Res_cascade[6];
assign Res_configs[8][3] = Res_cas_in_temp[4];
assign Res_configs[9][3] = Res_cascade[8];
assign Res_configs[10][3] = Res_cas_in_temp[5];
assign Res_configs[11][3] = Res_cascade[10];
assign Res_configs[12][3] = Res_cas_in_temp[6];
assign Res_configs[13][3] = Res_cascade[12];
assign Res_configs[14][3] = Res_cas_in_temp[7];
assign Res_configs[15][3] = Res_cascade[14];
assign Res_configs[16][3] = Res_cas_in_temp[8];
assign Res_configs[17][3] = Res_cascade[16];
assign Res_configs[18][3] = Res_cas_in_temp[9];
assign Res_configs[19][3] = Res_cascade[18];
assign Res_configs[20][3] = Res_cas_in_temp[10];
assign Res_configs[21][3] = Res_cascade[20];
assign Res_configs[22][3] = Res_cas_in_temp[11];
assign Res_configs[23][3] = Res_cascade[22];
assign Res_configs[24][3] = Res_cas_in_temp[12];
assign Res_configs[25][3] = Res_cascade[24];
assign Res_configs[26][3] = Res_cas_in_temp[13];
assign Res_configs[27][3] = Res_cascade[26];
assign Res_configs[28][3] = Res_cas_in_temp[14];
assign Res_configs[29][3] = Res_cascade[28];
assign Res_configs[30][3] = Res_cas_in_temp[15];
assign Res_configs[31][3] = Res_cascade[30];
assign Res_out_temp[0][3] = Res_cascade[2];
assign Res_out_temp[1][3] = Res_cascade[4];
assign Res_out_temp[2][3] = Res_cascade[6];
assign Res_out_temp[3][3] = Res_cascade[8];
assign Res_out_temp[4][3] = Res_cascade[10];
assign Res_out_temp[5][3] = Res_cascade[12];
assign Res_out_temp[6][3] = Res_cascade[14];
assign Res_out_temp[7][3] = Res_cascade[16];
assign Res_out_temp[8][3] = Res_cascade[18];
assign Res_out_temp[9][3] = Res_cascade[20];
assign Res_out_temp[10][3] = Res_cascade[22];
assign Res_out_temp[11][3] = Res_cascade[24];
assign Res_out_temp[12][3] = Res_cascade[26];
assign Res_out_temp[13][3] = Res_cascade[28];
assign Res_out_temp[14][3] = Res_cascade[30];
assign Res_out_temp[15][3] = Res_cascade[32];
//////////////
//conf_2
assign I_configs[0][2] = I_in_temp[0];
assign I_configs[1][2] = I_in_temp[1];
assign I_configs[2][2] = I_in_temp[2];
assign I_configs[3][2] = I_in_temp[3];
assign I_configs[4][2] = I_in_temp[0];
assign I_configs[5][2] = I_in_temp[1];
assign I_configs[6][2] = I_in_temp[2];
assign I_configs[7][2] = I_in_temp[3];
assign I_configs[8][2] = I_in_temp[0];
assign I_configs[9][2] = I_in_temp[1];
assign I_configs[10][2] = I_in_temp[2];
assign I_configs[11][2] = I_in_temp[3];
assign I_configs[12][2] = I_in_temp[0];
assign I_configs[13][2] = I_in_temp[1];
assign I_configs[14][2] = I_in_temp[2];
assign I_configs[15][2] = I_in_temp[3];
assign I_configs[16][2] = I_in_temp[0];
assign I_configs[17][2] = I_in_temp[1];
assign I_configs[18][2] = I_in_temp[2];
assign I_configs[19][2] = I_in_temp[3];
assign I_configs[20][2] = I_in_temp[0];
assign I_configs[21][2] = I_in_temp[1];
assign I_configs[22][2] = I_in_temp[2];
assign I_configs[23][2] = I_in_temp[3];
assign I_configs[24][2] = I_in_temp[0];
assign I_configs[25][2] = I_in_temp[1];
assign I_configs[26][2] = I_in_temp[2];
assign I_configs[27][2] = I_in_temp[3];
assign I_configs[28][2] = I_in_temp[0];
assign I_configs[29][2] = I_in_temp[1];
assign I_configs[30][2] = I_in_temp[2];
assign I_configs[31][2] = I_in_temp[3];
assign Res_configs[0][2] = Res_cas_in_temp[0];
assign Res_configs[1][2] = Res_cascade[0];
assign Res_configs[2][2] = Res_cas_in_temp[1];
assign Res_configs[3][2] = Res_cascade[2];
assign Res_configs[4][2] = Res_cas_in_temp[2];
assign Res_configs[5][2] = Res_cascade[4];
assign Res_configs[6][2] = Res_cas_in_temp[3];
assign Res_configs[7][2] = Res_cascade[6];
assign Res_configs[8][2] = Res_cas_in_temp[4];
assign Res_configs[9][2] = Res_cascade[8];
assign Res_configs[10][2] = Res_cas_in_temp[5];
assign Res_configs[11][2] = Res_cascade[10];
assign Res_configs[12][2] = Res_cas_in_temp[6];
assign Res_configs[13][2] = Res_cascade[12];
assign Res_configs[14][2] = Res_cas_in_temp[7];
assign Res_configs[15][2] = Res_cascade[14];
assign Res_configs[16][2] = Res_cas_in_temp[8];
assign Res_configs[17][2] = Res_cascade[16];
assign Res_configs[18][2] = Res_cas_in_temp[9];
assign Res_configs[19][2] = Res_cascade[18];
assign Res_configs[20][2] = Res_cas_in_temp[10];
assign Res_configs[21][2] = Res_cascade[20];
assign Res_configs[22][2] = Res_cas_in_temp[11];
assign Res_configs[23][2] = Res_cascade[22];
assign Res_configs[24][2] = Res_cas_in_temp[12];
assign Res_configs[25][2] = Res_cascade[24];
assign Res_configs[26][2] = Res_cas_in_temp[13];
assign Res_configs[27][2] = Res_cascade[26];
assign Res_configs[28][2] = Res_cas_in_temp[14];
assign Res_configs[29][2] = Res_cascade[28];
assign Res_configs[30][2] = Res_cas_in_temp[15];
assign Res_configs[31][2] = Res_cascade[30];
assign Res_out_temp[0][2] = Res_cascade[2];
assign Res_out_temp[1][2] = Res_cascade[4];
assign Res_out_temp[2][2] = Res_cascade[6];
assign Res_out_temp[3][2] = Res_cascade[8];
assign Res_out_temp[4][2] = Res_cascade[10];
assign Res_out_temp[5][2] = Res_cascade[12];
assign Res_out_temp[6][2] = Res_cascade[14];
assign Res_out_temp[7][2] = Res_cascade[16];
assign Res_out_temp[8][2] = Res_cascade[18];
assign Res_out_temp[9][2] = Res_cascade[20];
assign Res_out_temp[10][2] = Res_cascade[22];
assign Res_out_temp[11][2] = Res_cascade[24];
assign Res_out_temp[12][2] = Res_cascade[26];
assign Res_out_temp[13][2] = Res_cascade[28];
assign Res_out_temp[14][2] = Res_cascade[30];
assign Res_out_temp[15][2] = Res_cascade[32];
