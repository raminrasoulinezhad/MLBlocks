module template (

	);
	
	///////// Parameters

	///////// IOs

	///////// internal signals

endmodule 
